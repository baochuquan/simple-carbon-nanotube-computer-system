`ifndef _SIGNALS

`define sel_A_DI	2'b00
`define sel_A_acc	2'b01
`define sel_A_pc	2'b10
`define sel_A_x		2'b11
`define sel_B_DI	3'b000
`define sel_B_nDI	3'b001
`define sel_B_nacc	3'b010
`define sel_B_C		3'b011
`define sel_B_zero	3'b100
`define sel_B_x		3'b101

`endif